library ieee;
use ieee.std_logic_114.all;


entity overflowdetecter is

port(
a.b:in std_logic_vector(1 downto 0);
c:in 


);

end overflowdetecter;